library ieee;
use ieee.std_logic_1164.all;


entity AND_9 is
	port (A,B,C,D,E,F,G,H,I : in std_logic; Y : out std_logic);
end AND_9;

architecture BHV of AND_9 is

begin
	Y <= A and B and C and D and E and F and G and H and I;
end BHV;